module decoder_6_64(
    input  wire [ 5:0] in,
    output wire [63:0] out
);

// 生成块
genvar i;
generate for (i=0; i<64; i=i+1) begin : gen_for_dec_6_64
    assign out[i] = (in == i);
end endgenerate

endmodule